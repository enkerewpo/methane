module midi.MidiProc(
  input   clock,
  input   reset
);
endmodule
