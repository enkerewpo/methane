module MidiProc(
  input   clock,
  input   reset
);
endmodule
